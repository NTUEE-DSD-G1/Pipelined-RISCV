module show;
    initial begin
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOkkkkkkkkkkkkkkxkkxlccccccccccccccc:::::::::::cloolloooooooooooooo");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOkkkkkkkkkkkkkkkkkkkxxxxxlcccccccccccccccccc::::::::coddoloollooooooolll");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOkkkkkkkkkkkkkkkkkkkxxxxxxxxocccccccccccccccccccc:::::cokkkkkkxoloooooollll");
        $display("OOOOOOOOOOOOOOOOOOkkkkkkkkkkkkkkkkkkkkkkxxxxxxxxxxxxxoccccccccccccccccccccccc::cloooolddolllllllllll");
        $display("kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkxxxxxxxxxxxxxxxdddolcccccccccccccccccccccc:ccllllc:oollllllllllll");
        $display("kkkkkkkkkkkkkkkkkkkkkkkkkkxxxxxxxxxxxxxxxxxxxddddddddolccccccccccccccccccccccccllllllodollllllllllll");
        $display("xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxdddddddddddddddddolccccccccccccccccccccccccllllllodlllllllllllll");
        $display("dddddddddddddddddddddddddddddddddddddddddddddddddooodollclccccccccccccccccccccclooooodollooooooooooo");
        $display("dddddddddddxxxxxxxxxxxxxxxxxxxxxxxxxddddddddddddddxxxxolllllllllllllllllccccccloooooodoloooooooooooo");
        $display("dxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxdxkOkkOkOkolllllllllllllllclccccccoodooloddooddddddddddd");
        $display("xxxxxxxxxxxxxxxkkkkkkkkkkkkkkkkkkkkkkkkkkkxkxkxddxxxxxdoooooooooooooooodooododxxxdoldxxddxxxxxxxxxxx");
        $display("xkkkkkkkkkkkkkkkkkkkkkkkkkkOOOOkkkkkkkkkkkkkkkxcokkkkkkxxxxxxxxxxxxxxxkOkxxxxxxxxoclxxkxdxkkkkkkkkkk");
        $display("kkkkkkkkkkOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOklokOkkkkkkkxxxxxxxxxxxxx00kxxddoccc:lxxkkxkkkkkkkkkkk");
        $display("kOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOxdkOOOkkkkk00Okxxkkkxxxx0XOxxxdl',lddxxxxdxkkkkkkkkkk");
        $display("kkkkkkkOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOkkkkkkkxxkkkxkxxOXNNX0kxddooook0koooll:coxdooollclooddddddd");
        $display("xxxxxxxxxxxxxxxxxxxxdxxxxxxkkkkkkkxxxxxxdoollc:cddoooolllx00KNNX0Okkxxxkxxxdddxddxkxxxoc:lxkkOOO0000");
        $display("dddddddddddddddddddoodddddddddddddddl:::;,''....'coc::::;lkxx0K0kkkkkkxxxxxxxxxxdxxxxdc;:odddddddxxd");
        $display("xxxxxxxxxxkkkkkkkkkxxxkkkkkkkkkkxxo:,'....    ....'''''',:oooooxxxdddodxkxdolllllllll:;;cloooooodxdd");
        $display("OOOOOOOOOOOOOO0000OOO00000000000x;...                  ...',::;:loolccclxxdolcccccclc;',:ccllclcllll");
        $display("OO00OOO0000OO00KKK000KKKKKKKKK0d'                         ...;ccccc::cc:cloolllllcllc,,cllllllllllll");
        $display("0000kk0KKK0kkKKKKKKKKKXKXXKK0x:.     ...''.......           .'loooolllllollcccclllooc;colllloooooooo");
        $display("OOOOOkOOOO0OO00000000KKKK0Oxc,'''....''',,,'''''''''...     ..,oddoollooddooolllllllllllllllllllllll");
        $display("0000O0000000000000000K000koc:c:;'...''..;:;,''...',,,,'..   ...:dkkxxxxxxxxxxxxxdddddddddddddddddddd");
        $display("XXXXXXNNNNNNNNNNWWNNWWNNNOcokd;..'....,col:,''..'',,',::;.   ..,oOKK0OOOkkkkkkxxxxxxxxxxxxxxdddddddd");
        $display("XNNNNNNNNNNNNNNNNNNNNWWNN0llkd:;;;;,,;:cllc;,,,,,;::c::col,.  .;lOKKKK00OOkkkkxxxxxxxxxxxxxxxddddddx");
        $display("XNNNNNNNNNNNNNNNNNNNNNNNWO,'odlcc:;,'.','.,::;;;;:::cldddxd;....;kXXXXKK000OOkkkxxxxxxxxxxxxxxxdl:::");
        $display("XNNNNNNNNNNNNNNNNNNNNNNNNk:clc::::;,..','..,;;;::ccclooxkkxl'.. .oKXXXXKKKK000OOOOOkkkkkkkkOOOkx:...");
        $display("XXNNNNNNNNNNNNNNNNNNNNNNNOl:;:::::;,,,,,;:cccc:;:cclooddxxxd;....;xKNNXXXXXXXXKKKKKKKKK0000Okkxdc;;c");
        $display("XXXNNNNNNNNNNNNNNNNNNNNNNOc;;;::::;'......':ooc::ccllooodxxd:.  .'okKNNNNXXXXXXXXXXXXXKKKKK00Oxdllod");
        $display("XXXXNNNNNNNNNNNNNNNNNNNNXx:;;;;;;,..''.''...':c:::cccllloddd:.   'dO0XNNNXXXXXXXXXXXXXXXXKKK0kxdoood");
        $display("XXXXNNNNNNNNNNNNNNNNNNNNKo:::;;,'.....'.......,;::c::::cllooc,...,kKXNNNNNXXXXXXXXXXKKKKKKKK0Okxxddd");
        $display("XXXNNNNNNNNNNNNNNNNNNNNN0l:::;,'.  .......   .';::cc:::::cllc:;,':ONNNNNNXXXXXXXXKK000OOOOOOkkkkxddd");
        $display("XXNNNNNNNNNNNNNNNNNNNNNN0l:::;,''. ..   ....',;;::::::::::cl:,;;,c0NNNNNXXXXXXXXXKK000OOOOkkkkkkkxdd");
        $display("XXNNNNNNNNNNNNNNNNNNNNNN0l:::;,,;,''....,:clllc::::;:::::::c:,;ccdXNNNNNNNXXXXXXKKKK000OOOOkkkkkkxdd");
        $display("XXXNNNNNNNNNNNNNNNNNNNNNOl::;;;;;;;;,,,;:cccccc::;;;;::;;;::coooxKNNNNNNNNXXXXXXXKKKK000OOOOOkkkkxxx");
        $display("XXXNNNNNNNNNNNNNNNNNNNNN0dl:;;;;,,,,,,,;;;::ccc::;;;;;;;;;;..:dkKNNNNNNNXXXXXXXXXXKKKK00OOOOOOkkkkxx");
        $display("XXXXNNNNNNNNNNNNNNNNNNNNNN0l;;;,,,,''''',,;:::::::;;;;;,,,. 'kXXNNNNNNNNXXXXXXXXXXKKK000OOOOOOOOOkkx");
        $display("dddxxxxkkO0000KKKKKKXXXXXXXkc;,,,''.....'',;:::::;;;;,,,,. ;0NNNNNNNNNNNNNNKOxxxddxO0OkOOkxddoollloo");
        $display("...''',,,,,::ccccccllloooolc;''.........',,,',,,,''''''''..cdooddxxxxxkkxddl,,;;;;;:;,''''.......,;;");
        $display("............'',,,,,,'''''''..............','..................................'.......    .......,,,");
        $display("...........................................'...............................             ........''..");
        $display("........................ ..............................................        ..............''...  ");
        $display(".................      .................................................    ...................     ");
        $display("............       ...............  .................. .....................................  ......");
        $display(".....           ................   ............................         ............................");
        $display("..........................'.....  ....   ....  ..............       ................................");
        $display("  ................. .........   ........    ..    ........        ..........  ......................");
        $display("  .............. .   .....        .......  .............       .............    ....................");
        $display(".................. .....          ....................        .............     ....................");
        $display(".....   ......    ...            ......  ............       ...............     ...;;'..............");
        $display("\n\n\n");

        $display("MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM");
        $display("MMMWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWMMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWWWWWWWWWWWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWWWWWWWWWWWWWWWWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWNNWWWWNKOkkxdoolllodxxkOKXNWWWNNNNWNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWWNKko:,...............',;cdk0XNNWWNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNXOoc,.........................':d0NWWNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN0o;...............................';dKNNNNNNWWWNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKo,....................................;d0NNNNWNWWNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNXx;.......................'................,ckXNNWWWNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNXo'....................,;cclllllllllllllc;.....cONWWNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNXo....................;lxkOOOOOOkkkOOOOOkxxo,....'dXNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNx'..................,lxO00000KKKK000K0000OOkx:.....oXNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNO;.................';okO000KKKKXXKKKKKKK0000OOx;....'xNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNKc................,codkOO00KKKXXXXXXXXXXKKK0000Oo'....:KWNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNk,.............,:ldkkkOO00KKKXXXXXXXXXXXKKKK0000x:....;0WNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNd'..........';lodxkOOOOO00KKKXXXXXXNNXXXKKKKKK00Oc....;0WNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNXo..........,:lddxkkOOO000KKKXXXXXXXNNNXXKKKKKK00Oo'.'.cKWNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNXl.........,:lodddddddxkkO0KXXXXNNNNNNNNNXXKK00000d'.';kNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNXo..'......,codddoooddxxxxxkO0KXXXXXXXXK00OkkkkkOOd..'oXNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNk:,,,'....,:cclodxO00000OOOO000KXXXXK0O0000KK0OkOd..:ONNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNKxcll,...':oooodk00OkkdllxkkOkdxO00kkOOxdxO0kOOOkl',kNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNOddo:...,codxkkO00OOOkxxOOOOdloOXOdx00kddOOxkO0OdcxXNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNW0xdoc;',:lodxkOO00K00KKKK00Okxk0XKOO0KKKKKKK0000doKWNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNWNOxxdc:clldxkOO0KKKKKKKKKK0OOOOKXXKKKKKKKKKKKK0KOOXNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNWXOkkolllodxkO0KKXXXXXXXXK0OkO0KXXXXXXXXXXXXXXKKKXNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNWWXOkdloooddxO0KKXXXXXXX0kOOkO0KXXXKKKKKXXXXXXKKXNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWNkcloooddxxkO0KXXXXXK0kdkOOO0KXXKKKKKK0KXXXKKKNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWk.'ooodxkkkO0KKKKKKK0OkkxkkkO0K000KKKKKKKKKKXNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWXd:ldddxkOO00KKKKK00OO000KKKKKXXKKKKKKKKKK00XNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNWNNWN0doddxkO00KKK000kdxkkOOOOO000OOOO00KKKK00KNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNWN0l;coodxkOO0KKKKKOdoxO0KKKKXXK0kodO0KKKK0KNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNXOo:',colodxkkO000000OxdxkOKK0000OkOKXKKK00KXNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNNNNNNKOkdl;,,';odlllodxkO00000OOkxkkOOO0OOO0KKKK000KNNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNNNNNNK0kdl:;;,,,,,,:dkxolllodxkO00OO00OOOOOOO00KKKKK00KXNNNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNNNNNNX0kxoc:;;,,;;,,,,,,cxOOkxooooddkOOO00KKKKKKKKKXXKK0kxO0XNNNNNNNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNNNNNNX0Oxdlc:;;:;;;;::;;,,,,;cx00OOkxdooodddxkO0KXXXXXXXXXK0xoooooxkO0KXNNNNNNNNNNNNNNNNNWMM");
        $display("MMWNNNNNK0Oxdlcc::::::::::;::::;;,;;:cxKK00K0OxdddddddxxkO0KKKKK0OKkllooooolllodkkO0KXNNNNNNNNNNNWMM");
        $display("MMWXKOxdllc:cc:cccccc::::;,:::::;;;;:cd0K00KXXK0OkxxxxxxxxxkOOkO0KXkllooooolllloolloodxO0XNNNNNNNWMM");
        $display("MW0oc::cccc::c::ccccc::::,;:cc:::;;;:coO000KKXXXXKK0OkkkkOOOO0KXNNNKdlooolllllllllllllllldk0XNNNNWMM");
        $display("MWk::cc::::cc:::cccccccc:;:ccc:c:;,;::o0XKKKKKXXNNNNNX0OkkOKXNNNNNNNklooollloolllllllllllllldkOKXWMM");
        $display("MWk:::::cccccccccccccccc::ccccccc::;::ckXNXXK0KKXNNNNNNKkOXWWNNNNNNN0olollloloolllllllllcccclllld0WM");
        $display("MWk:::::::::cccc::ccccc:;:lccccllc:;:cco0NNNNXKKKXXNNWXOxxkKNNNNNNNNKdlollloollllllllllllllccllcckWM");
        $display("MWk:::::::ccccccccccccc;;ccccccclc:::cccoKNNNNNXXKKXX0ddxdll0NNNNNNNXxcolllllllllllllllllllcccccckWM");
        $display("MWk::::::::ccccccccccc:;clcccccccccccccllxNNNNNNXXXX0c':dd::dKNNNNNNXxlllcccllllllllllccccccccccckWM");
        $display("MWk::ccc:cccccccccccc:,:lcccccccccccccccco0NNNNXXXXK0d;'locdkOXNNNNNXxclcccclllllllllccccc:cc:ccckWM");
        $display("MWk::cc:::cccc:::ccc:;,;cccccllccccccc:cclxXNNNNXKKKKd,'clckKK0XNNNNNkccllccclllcclcccccclcc::ccckWM");
        $display("MWk:::::::ccc::::ccc:c:;,;;cccccccccccccclo0NNNNXKKKk;.,cloxKNKKXNNXXkcccccccccccccc::cccc:::::::kWM");
        $display("MWkc:::::::c::c:c:::::ccc;,';ccccclllcc:cclkKXNNX00x;..,coodONNXKXXNXxcccc::cc::c::::::::::::::::kWM");
        $display("MWk:::;:::c::::::::c:::::;,;:cccclccccc:cclxOKNNKxl;'.';clood0NNNXXNXkc:c:::::::::::::::::::::;;:xWM");
        $display("MWx;::;::::c:::c:::::::;,;:cccc:cccccc:ccccdkKNXk:,,'',clodocxXNNNXXXx::c::::::::::::;::::::::;;;xWM");
        $display("MWx;;:;;;::cc::c::::::;,;cccccc::ccccc::cccld0NKl,,''';coddocl0NNNXXXk::c::::::::::::;;:::;:;;::;xWM");
        $display("MWd',;;,,;:cc::::::::,';::cc::::cccc::::cccclOXkc,,'',;clddolckXNXXXXk:;::::::::::::::;::;;;;;;;;xWM");
        $display("MWd...';,';::::::::::,.':cc::::::c::::cccccclOKo:;,'',;:lddoocdXNXXXXx:;::;:::::;;;;;:;;;;:;;;;;,dWM");
        $display("MWx'....'..,;::::::::;'.,:cccc::::::::cc::::lOkc:;,,,,;:looooloKNXXXXk;;::;;;;:;;,,;;::;;;;,;;,,,dWM");
        $display("MWx,''......';:;::::;;,..;:::::::::cc::cc:::cxdcc:;;;;;:looddoo0NXXXX0c;:::;;;::;;;,;;;;;;;;;;;,,dWM");
        $display("MWx;,,,''.. ..,;;::::;;,..;::::::::c::c::;;::odlc:;;;;;clooodooONXXXXKl,:::;;;::;;;;;;;;;;;,,,;,'dWM");
        $display("MWx;,,,,,''.  .',;::;;;;'.';::::::::::::::::ccllc:::::::looodooOXXXXXKl,;:;;;;;:;;;;;;,;;;;;;;,''dWM");
        $display("MWd',;;;;,,'.. ..,;;::;;,..';::c::::::::::::c:clc::::::clooooooOXXXXX0o,;;;;;;;;;;;;;;,;;;;;;,,''dWM");
        $display("MWo.',;;;;;;,'.  .,;;;;;;,..;:::::::::cccc::::clccc:c::cllloddokXXXXK0o,,;;;;;;;,;;;;,,,;;;;;,,,,xWM");
        $display("MWo..,,;;;;;;;;,...,;::;;;,..;;::cc::::::::::cccccccccccllloddoxKXXXKOo;,::;,;;;;;;;;,,;;;;;,,'',xWM");
        $display("MWKkkOO000000000OkkO0000000OkO0000000000000000000000000KKKKKKKKXWWWWNNK0O000OO000000OOO00000OOkkkKWM");
        $display("MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM");
        $display("\n\n\n");

        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO000000000000");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO000000000000000000KKK");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO000000000000000000000KKK");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO00000000000000000000000KKKKK");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO0000000000000000000000KKKXXX");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO0000000000000000000000000000KKKKXXNN");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO0OOOOOOOO0000000000000000000000000000KKXXNNNN");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO0OOOO00000000000000000000000000000000KXXNNNNN");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO00O0OOO000O0000000000000000000000000000000000000000KKXXNNNNN");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOO00O00000O000OOOOOOO000000000000000000000000000000000000KKKXXNNNN");
        $display("OOOOOOOOOOOOOOOOOOOOOO000000000000OOOOOOkkxxxxxxddddxxxdxkOO000000000000000000000000000O0000KKXXNNNN");
        $display("OOOOOOOOOOOOOOOOOOOOO00000000000OOOkkxdodddoooooooooddlccloxkkkOOO0000000000000000000OOOO0KKKKKXXXXX");
        $display("OOOOOkkkOOOOOOOOOOO00000000000OOkkkxdoddollollooolcc::ccclooodoodxkkO00000000000000000000XXXKKKKKKKK");
        $display("OOOOOkOOOOOOOOOOOO00000000000OOkddddddolccll:cc:;,,,:lolcllcccclclodxO000000000000000000KKXK0KKKKKK0");
        $display("OOOkkOOOOOOOOOOOO000000000OOOkxlccccc:;,,,;,',,,'',,:cc:::,,:lllllcloxkO0000000000000000000000000000");
        $display("OOkkOOOOOOOO000000000000OOkxol:;;,',,''''''''''.'',,,,,,,'',:clcclooodxkO0000000000000000000OO000000");
        $display("OkkOOOOOOO000000000000Oxdool;,,,''''...''.......'''....''',,;;;,:loddoxOOO00000000000000000OxdO00000");
        $display("kOOOOOO0000000000000Oxoolc:,'','.'......................'''''''',:clocokO0000000000000000000OkxO0000");
        $display("kOOO000000000000000kdllc:;'..'.................................'.,::c::oxO0KK00000000000000000kxk000");
        $display("OO000000000000000Oxl:c:'''.......................................',,:;;cldxOKK0000000000000000OkxkO0");
        $display("O000000000000000ko:;;;'..........................................''',,,;:llokO0KK0000000000000OOkxxO");
        $display("000000000000000Oxl,,,..............................................'''',:cccooxO0O000000000000OOOOxx");
        $display("O00000000000000kdc,''......................................'''.......''',::::clxkOO00000000OOOOOOOOx");
        $display("000000000000000ko;'''.....................................',,''..''.''..',;,;;:okO00000000OOOOOOOOOO");
        $display("OO00KKK0000KK00kc'.'....................................',;;;,,'''''''..',,''';lxO00O000OOOOOOOOOOOO");
        $display("OOOOO00KKKKKKK0kc.......,'....'.............''........',,;:::;,'''',,''',,'..',lkOOOOOOOOOOOOOOOOOOO");
        $display("OOO0000000KKKK0kc'....,;::;,',,'',,,'''...',,,''.....,;;;::::;,'.',;;,,,;;'..':xOOOOOOOOOOOOOOO00000");
        $display("OOOOO0000000000kl,...';cclc:;;,,'',,''''',,;:;;;,'.';:::;::;,,'..',,;:::::,'';lk0OOOOOOOOO000000000K");
        $display("OOOOOOO000KK000ko,'..'clllc::;;;;;;,,'',,,;::::c:,,,:::;,,,,,,'',;;;::ccc:,,,:okOOOOOO000000000KKKKK");
        $display("0000OOOOOO00KKKKx:,'',;:ccclloooooollcccccc:::clc::;;;::::cclccclllllllool:;,;lk00000000000KKKKKKXXX");
        $display("000KK0000OOO000K0xc,,;:cooodddddddoolllllool::::::;;;:clllllllllllllllloollc;cx0000000KKKKKKKKXXXXXX");
        $display("KKKKKKKKKKK000O000ko:c:codoolc:cl:;,,:ccclolc:cllcc:::ccc::;,,,;c:,;:cloddOxlkK00KKKKKKKKXXXXXXXXXXX");
        $display("KKKXKKXXXXXXXXKK000kloxoddolc::cc:,,,;::cllc::looolc::ccc::;,,,;ccccclodxk0ko0KKKKKKXXXXXXXXXXXXXXXX");
        $display("XXXXXXXXXXXNNNNNNXX0olxxxddooooooolccclllllc:cooddooc:;clllllcllooodddxxkOOdxKXXXXXXXXXXXXXXXXXKKK00");
        $display("NNNNNNNNNNNNNNNNNNNXdcoxxxddddddddoooooooolccoodddddoc:coooooloooodddxxxkOdlkKXXXXXXXXXXXXKKKK00000O");
        $display("NNNNNNNNNNNNNNNNNNNXKkddxxddddddddooooddoolloodddxxddolclooooooodddddddxxddk0XXXXXXXXKKK00000OOOkkkx");
        $display("0KKXXNNNNNNNNNNNNNNNNXOdddxxxxddddddddoolloooddxxxxxxdollcllooooddddddooodkKXXXXKK00000OOOOkxxxxkOO0");
        $display("OOO00KKXXXNNNNNNNNNNNNKkddoddooooooooolllllodddxxxxxxxdolccllllooooooooodxOKK00000OOOkkxxxxkkOOOO0XX");
        $display("OOOOO0000KKXXXXNNNNNNNX0xxxddddoooooooooloodddddxxxxxxxxdolloodddddddddddxO00OOOkxxdxxkkOOOkxkOOOOKX");
        $display("OOOO000000000KKKXXXNNNNKkxxxxxdddddddoolodddooddddddddooddollooddddddddddxkOkxxxkkkOO00OOkOOkOOOOxod");
        $display("OOOOO0000000000000KKKXXX0xxxxxxxxdddddoooolc::llooollc;;cllooodddddddddodxkOOO00kkOOkkkkkkxdllooddc:");
        $display("OOOOOOOO00000000000000000kddxxxdddddddddooollooooooooolllooddddddddddooox0000OOOO00Oxdlc;::,;:cloxkx");
        $display("O00000OOOOOOOOOOO00000000OxddxxxxxdddddddddoodddooddooddddddddddddoooolodddxkOOxdl:;'...,:odxxkkOOOk");
        $display("O00000000000OOOOOOOOOOOOOOkxddxdxxxdddddddddddddoddddddddxxxddddooooolokkkOkdoollc:cclldddx00O0Oxddo");
        $display("000000000000000OOOOOOOOOOOOkxdddxxxdddddddddddddddddddddddddddddooolloxOOkO0OolxxdddddoolccxK0K0dlll");
        $display("O0000000000000000000OOOOOOkkxdddddxddddodddoolllllllclloooooloooolllodxO0kxxkxxdollccc:;;;';O00XOoll");
        $display("00OOOOOO0000000000000OOOOOOkxxddddddddooolcc::::c:::;;;;::cccclllllldOOxooolccc:::;;,''';:,'oK0KKxll");
        $display("0000kxkO00KKK00000000OOOOOOOkkxddddddooll:;;;;;;::::;;;;;;:::cllllloxkxdccol:,',,,,,,..,loc,;O00X0dl");
        $display("odxOkk00000KKKKKKK0000000OOOOkkxxdddddooolcccccccccccccccccccllllloodxxxdlllolcloollc:;:odol:dK0KKkx");
        $display("co0XKKKXXXKKKXXXKKKKKKK00000OOOkddddddddooolllccc::cccccccccllllllllodxl;:::cc::clooooooxxxkxx000KKk");
        $display("okKKKKXXXK000OKXXXXXXKKKKKK00Okdoc:lddddoooollllcccccccllllllllllcccldo:,,',;,'',,;;::ccloddxxkOkO0k");
        $display("xkOO0KXXKOxxxxO00KXKKXXK00Oxolloc'.'coooooooolllcccccccclllllclc:::::c:,'..'......'',,;::cclllloddxx");
        $display("xkkkKNXNXkoxkOkxxxxxkkxdoddo:,:lc'. .cooooololllcccccccccllccc:;;:;;;,..............',,,;;;;;::clood");
        $display("dkxkO0KXKkxkO0Oxxdolc:;;:cll:,;cl;. .'cooolllllccccccc:cclllc;;;,,,;'.............''',,,,,''',,,;;:c");
        $display("xdoooloxK0xodolcccc:;'',,,,;,,,;cc,..',:llllllccc::::::cccc;,,;,''...................'''''''''''''''");
        $display("odddodkO0Odc::;::::;,,'''',;,,'';c:;;;'';:ccccc:::::::::;;,,;;,'.....  ......''..........''........'");
        $display(":lllokOOxl:;;;;;::;,''.',,,,,,'..;c:;;,..,;::::::;;,'',',',,,'....    ............................',");
        $display(";;',:loo:;,,;,,,''.....'',''''....''.,;'..',,,,,''.''''',,'.....     .........................'''',,");
        $display(":;';clc;,,,,,',;,...''''''''''.........'......'''...',,,''.        ...........................''''',");
        $display(":;,;:c:,,,,,,,;;'..'''''''''.........................','..       .................................''");
        $display("'....,,,','',,,,'..''...''...................  ... .....       .....................................");
        $display(";,,',,''.''',,,''...'........................               ........................................");
        $display("ooolc,.....',,'''..''.........................          ............................................");
        $display("dodo:'.....,,'''...''.........................  ..  ................................................");
        $display("dddo,.'...',,''..'''................................................................................");
        $display("xxdc,'....'''''''...................................................................................");
        $display("xxo:,'....'''''''...................................................................................");
        $display("\n\n\n");

        $display(",,;;;,;;,,,,'.......'::;;,.',,,,,,,'.........;:;;;;;;cccccccllcccccccc:,''''''''''''''''''''''''''''");
        $display(";;;:;;;;;;;;'.......;::;:c:c;,,;;;;,........'::;;;:::clcccccclccccccclc,,,,'',,'',,,,,,,,,,,,,,,,,,,");
        $display(":::::;;:::;;,......,::ccc:cc;;;;;;;,........';;,,;;::llccllloollllolooc;;;;;,,,,,,;;;;,,,;;;;;;,,,,,");
        $display("::;:c:::::::;......,:,,::;:c:;;;:::,.................,:cllooddddddddddc;;;;;;;;;;;::::;;;;;;,,,,,,,,");
        $display(";,,';l::::::;......;:;;c:;clc::cccc;..'::;',,'....... .;oodxxkOOOkkkkdc:::::::;:::::::;;;;;,,,,,,,,,");
        $display(",,''ldc:cc::;'.....,c;;cc:lolclllll;'':ol;',;'....'.''':oddxkkOOOkkkOdc::::::::::cc::::;;::;;;;,,,;;");
        $display(",,,;dxolllllc,.....,c::llcodooooddo;...,:c::,'......,ldxxxkkkkOOkkkkko:::cclcccccccc:::::c::::::::::");
        $display(":::cO0dooollc,.....;lllooodddddxdddl:ccc:;:;,'''''''';::ccclloddxxxkxocccclollollllllccccccc::::cc::");
        $display("ccclOKkdddooo;''''';lolcldkxddxddddddxxolllc;;;:::;;::::c:::::cc::coolccclooolllloollccc::cccccccccc");
        $display("looo0X0kkxxdo:''''':oododkOkocldxkkxxxdoolllloddoooollccc:c:;:::::::cccllolllllllllcc:::ccccc::cc:::");
        $display("oodd0N0Okkkxxc,,,,,cxkkddxxdoc:lxxddlloolclodxdlloddolc:::;,,:cccccc:clcccclooollolllcccllcccclc::::");
        $display("ddxx0NKOOOkkkl;,,,,lxkxxdoc::;,:lddoloodllddxdlcllooooc::;;,',:cllc::cccccllooooooooooollccccclllllc");
        $display("kxxx0NXK0OOOkdlcccclxkOOkl:,'';lxxdoooooddxxdolclllloooc::;,'.';::;'':oooodddoooooooooollllllllllllc");
        $display("OOOOKXXK0000OOOOOOOkkkkkxoc;,';xkxdddxxkxddooollllllllllc:;,'.,;;,',:oddddddddddollllllcccclccccc:::");
        $display("KKKKK0000000000OOOO00OOOkxoc;''cdxxxkkkkxooolllllllllccccc:;,;:;,,cddddodddoodoolllcclllccccccccc:::");
        $display("0000000OOOOkOOOOOOOOOOOkkkkxl;,,;cloxkkkxddollllllllcccc::;::;,,;lolcloddddddoooooooddoolllllllllccc");
        $display("OOOOO00000OOOkkkkkkkkkkkkOOOkdl:;,'.',,,,,,,,,'''''',,,;:;;,,'':xx:...:ooodoododoooodooooooooolcccc:");
        $display("000000000OOOOOOOOOOOOOkOkkkkkOxc,'.......   ..      ..',,,'....;xd:,''coooooddodddoooolloooooollcc::");
        $display("KKK0000000000000000000KKK0000OOxc'.......   ....... ........  .cxxdddddxddddddoooooooolllloooolllccl");
        $display("KKKKKKKKKKKKKK000KK000000000000K0d;....     ..........       .;xkxxdxxxxddxdddooooooollllooooooollll");
        $display("KK0KKK000KKKK0000000000000000OOO0Oo;'.......;c,........     ..lkkxxxxxxxxxxddddddddooooolllloollcc::");
        $display("0000000000000000OOOOOOOOO000000OOOOxl;''''..:kkdolll;''......,ldddddxxxxxxddddddddddddolllllllllcccc");
        $display("OOOOOO00OOOO00OOOOOOOOOOOOOOOOOOOOOOxc,,''':xOOOOOOOdc::;;''.'lollcccccllloooddddoooooollllllllllllc");
        $display("OOOOOOOOOOOOOOOOOOOOOOOOOOOOkOkkOOkkxolc:;,;dkkkkkkkkdc::;,.'cxxxddoollcc:::::ccllllloolollllccccccc");
        $display("kkkkkkkkkkkkkkkkkkkkkkxkkkkxxxollc;'........,clooooooooxdl:,;looooooooooollcc:::;;;,,,;;::::ccccccc:");
        $display("xxxxxxxxddxxxxxxxxxxxxxxxxdl;.........'',;;;:::ccccccc:cc;,..';;::::cccccccccccccc::;;,,'''.''',,,;;");
        $display("oooodddddoddoddddddddddddddollcccclllloooooooooooooooo;.      ...',;;;:::::::::c:::::ccc:;;;;;,'','.");
        $display("llllllllooooooooooooooodooodddddddooooooooooolooollllll:.....   ..',,;:::cccc::::::ccldxoododxdoddc,");
        $display("\n\n\n");

        $display("00000000000000000000000000000000000000000000000000OdlodxxkO00KKKKKK00000OkkkkkOO0KKXK000000000000000");
        $display("000000000000000000000000000000000000000000000000000kllddxkkO00KKKKK0K00OOkkkkkO00KKXK000000000000000");
        $display("00000000000000000000000000000000000000000000000000KOoloddxkO00KKKKKKKK0OOkkkkOO0KKKKK000000000000000");
        $display("0000000000000000000000000000000000000000000000000000xlloddxkO00KKKKKKK0OOkkkOO00KKKK0000000000000000");
        $display("OOOOOOOOOOOOOOOOOOOOOOOO0000O000000000000000Oxddxdooc:;:;;:cldk0KKKKK00OOOkOOO00KKK00000000000000000");
        $display("OkddxkOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOOkxdollc;'.'''............,cdk0KK00OOOOOO00KKK0OOOOOOOOOOOOOOOOO");
        $display("KklldkOkkkOOOOOOkkkkkkkkOOkkkOkkkkxdoc:,'........................';ldkOOOOO000KKK0OOkkkkkkkkkkkkkkkk");
        $display("NKOOOO0OOOOOOOOOOOOOOOOOOOOOOOkxoc;,'''..............................';codkO0KKKK0Okkkkkkkkkkkkkkkkk");
        $display("NKOO0XXXXXXNNXXXXXXXXXXXXXXK0xl;''..'...'................................';cdk000OOOOOOOOkkkkkkkkkkk");
        $display("dllodkO0KXNNNNNNNNNNNNNNNNKx:''........''...................................';lx0XXXKXKKKKKKKKKKKKKK");
        $display("......',:cldk0XXNNNNNNNNXk:..................................'''..............',lOKXXXXXXXXXXXXXXXXX");
        $display(". ...........;lxkKNNNNXOc'..................................''.'''.....''.''...'',lOXXXXXXXXXXXXXXNN");
        $display("     ..  ......',cxKNKo'........  ......    ........ ............''....',''''..',,,;d0XXXXXXXXNNNNNN");
        $display("   . ... .  ......'co;.................         .... .    ..............',''''..',,,;lOXXXXXNNNNWWWW");
        $display("'....''.......  ....................            ......   .......................'',,,,ckXNNNWWWWWWWW");
        $display("ccccccc;,'..... .........  .........        ......................................',,',ckNWWWWWWWWWW");
        $display("oddxxddol:;;,,...........  ..........    .......................'''................'''',:kNWWWWWWWWW");
        $display("xkkkkkkkkddooc;....................... .............''''.......,:;,''.....'........''''''c0WMMMMWMMM");
        $display("kkkkkOOOOOOkko,... ...........................'','.',;;;'..''.,clc;;,,''',;'''......'..'',oXMMMMMMMM");
        $display("kkOOOOO000OOx:.... ..  ....................'',,;;,',:cc:;',,,,:odlcc:;,,,::;'''.........'':OWWWWWWWW");
        $display("ddodddxkkOOOo'...  ..   ..................',;:::;;,;cllc:;;;;;ldxdollc:::clc;'''''..'..'.';oO00KKKKK");
        $display("cccloodxxxxd:....  ...    ...........''...,:cclc:::cooolllc:;cdddooollcc:cldc,'.'''''.','',lk00000OO");
        $display("lllodxkOOOOd;....  ..        .............,:loolccclddooddl:;:cllccllllccclddc'...'''.',,,;oKWWWWWWW");
        $display("lllcloxxO0Oo,..... ..       ..............';cooollodxxxxdoc::clodooddxddooooxdl;'''''.',,,;dXMMMMMMM");
        $display("looloxO00Oxc'.....         ....'''',;;,'...':lllooodkkkxdollloooollooodddxxxxkxo:,',''''',;xNMMMMMMM");
        $display("dddodxk0K0ko,....        ....''''',,;;;,''',;:clodxkOOkxolccc::::ccloooooddddxxxo:,',''',,:kWMMMMMMM");
        $display("ddddddxkkOOx;.....      ..'',,,,;;;;::cc::;;,,,;:cllllc:cclollc:::clooodxkOOxolxxo;'''.,,;oXMMMMMMMM");
        $display("ooodddxxkO0k:...........,;''''',,'..',;::cc:;,..';;;;,,lkxxdol:'..,cddccldxkko;:cxx:'''',:kNMMMMMMMM");
        $display("oloddxxkO00k;.....,xk, 'c;'''',::;'.';c::cc::,';ldxxxo:okkxxdoc:;;coddoodddddc,,;oOo,',,,lOXWWWMMMMM");
        $display("occlodxkOOOkc.....l0d'.,l:;,,;::cccccllllll:;',codxkOkoldxxxxdoooodddddxxxkkd:lxxoc,.',,:dOKXWMMMMMM");
        $display("olcclodxxkOkl'....':,',;::::::ccllllllllcc:,,,:loxxkOOkxooddxddodddxxxxxxkxdlokOOkc'':c::oO0KNWMMMMM");
        $display("ddolloddxxkx:.... .':;,,,,;;:::cccccccc:::;;;:codxkkOOOOkkxxdddddddddxxxkkkkO000Oxc,cxko:oO00KWMMMMM");
        $display("xddddddxxxxx:.......:c;;;;;::cccclllllllc:;::codxkkO0000OOOOkkkkkkkOO00000000000Od:cxOkocdO000XWWWWW");
        $display("clodxxxxxxkxc'......:l:;:::cclooddddoolc:::cccodxkkO00O00OOOOOkkOOO0000KKKK0000OkdcoxxxolxOO000KKKKK");
        $display("::codxxxxxkkl,''''.'cdc;::cclloodddoollc;:cc;',:oxxkxl:cdO0OOkkkOOO00000KKKK000OkxdxxxdodkOOOO000000");
        $display("dooddoddxxxkd;''''''lkl:;::ccloodddoolc:,;c:,.',coodxl,,:dkOOOOOOO0000000000000OkkxxxxdokOOOOOO00000");
        $display("odddoooddxxxxo;',,''lko:;;::cllooddddollc:c::cloddodxkkxdxkOOOOOOOO000000000000OOkOkkddkOkkkkOOO0000");
        $display("ooooooodddddxdl;'',,cxo:;;;:ccllooddoolllllcclodxxddxkkkkOO000OOOOOO00000000000OO0K0OkOOkkkkkOOOO000");
        $display("oooooooooodddxxxl;,,cdo:;;;::ccclloollccccccclodxdoodxkkkOOOO00OOOOOOOOOOOOO000OkO0000OkxxkkkkOOOO00");
        $display("llloooloooooddx0Kxl:cdd:;;;;:::ccccc::::::ccclldddoodxkkkOOOOkkkkkkOOOOOOOOOO00koodxxxxxxxkkkkkkOO00");
        $display("cccccclllloodxx0WNXKKKk:;;;;;::::::;;,,;;;;;:::clllooooodddxxxdddxxkkOOOOOOOO0OocloddxxxxxkkkkkkkO0K");
        $display(";;;:::cccloodxx0NWWWMW0l,,,,;;::::::;,....',;;;;:ccccclllloooolcloxkkkkOOOOOOOo,,,;clodxxkkkkkkkkkOK");
        $display(",,,,;;:cloodxxxkO0KNWWNx:,,,;;;;::ccc:;,,,;::ccllooooodddxxxxxxxddxkkkkkOkkkkl'..  ...',:ccldxxkOOO0");
        $display("'',,;:clooddxxxxxxOXNWW0l,'',,,;;;::::;;;;;;:clloooooddxxxxxkkkkkkkkkkkkkkxxl. .          ...',cxOOO");
        $display(",;;::cllooddddxxxxONNNNOl;'.'',,,,;;:::;;;;;::cccccccloddxkkkkkOkkkkkkkkxxxx:. ..            ..,cxOO");
        $display(";:::ccllooooddxxxx0NNNKd::,'...'',,;;;::::cccllloooooddxxkkkkkkkOOkkkkxxddxxl,,,;,,;,.      ..',,cxk");
        $display("::::ccllooooddddoxO0KKkc;,,,;,...',,;;::cccllooddxxxkkkkkkOOOOOkkkkxxdddxxxxo;,;;,;cc.     ..'',,,:o");
        $display(":ccccllol:,'''......','....','''...',;::cclllooodxxxxkkOOOOOOOkkkxxddddxxxxxdc:c:;,;;.    ..'',',,,;");
        $display("cllllll:..                       ...',;::clllooddxxxxkkOOOOOOkkxdddddxxxxxxxdc,,;::;,.  ..'''''''',,");
        $display(",;;;:;..                           ...',;:clloooddxxxxkkkkkkxxdddddxxxkkkxxdol;'...;:....'''''',,'''");
        $display("  ..                               ......',;:clooooodxxxxxdddddddxxxxkkxxxdolc;'.....'..''''''',''''");
        $display("                                    .........',;:ccclooddddxxdxxxxxxxxxxddolc:;'......''''''''''''''");
        $display("                                     ..........,:ccllodxxxxxxxxxxxxxxxddolc::;,'....''''''''''''''''");
        $display("                                      .........,:cllooddxxxxxxxxxxddddolc:;,,'.....'''''''''''''''''");
        $display("                                       ........',:clloodddddddddddoolc::;,'...........'''''''''..'''");
        $display("       ...                              .......',;::clooodddoooollc::;,'..............''''''''....''");
        $display("      ........                          .......',;::cclloooollcc::;,''..............''''''''''......");
        $display("      .........                        ........',;;::cccllcc::;;;,'................''''''''.........");
        $display("         ......        ...              .. .....',,;;;;;:;;;;,,'...................''''''...........");
        $display("        ......        ....               .. ..'''''',,,,,,,,,'.....................''''.............");
        $display("         ...           ...               ..  ..''''''''''''.........................................");
        $display(".....     .             .                 .. .......................................................");
        $display("...........             .                   ........................................................");
        $display("............            .                   ...........   ...........................''.............");
        $display("..............          .                    .........      ........................................");
        $display("................                               .....          ....................................'.");
        $display("..................                              .....           ..'...............................'.");
        $display("\n\n\n");

    end

endmodule